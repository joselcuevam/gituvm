//////////////////////////////
//
//
// Comments here added
// branch1 done
//
/////////////////////////////
task testing_task;
 input a;
 input b; 
 begin

 end
endtask
//////////////////////////////
//
//
//  added a new message here
//  removed the previous one
//
/////////////////////////////
