//////////////////////////////
//
//
// Comments here added
//
//
/////////////////////////////


task testing_task;
 input a;
 input b; 
 begin

 end
endtask
