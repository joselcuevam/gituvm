
task print_message;

  input [7:0] a;
  input [7:0] b;
  
  begin

  end

endtask
